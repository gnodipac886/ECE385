module control(input logic clearA_loadB, );