module datapath ();

endmodule 