module ALU(
			input logic 	[15:0]	A, B, 
			input logic 	[1:0]	aluk,
			output logic 	[15:0] 	ans
		   );
	
endmodule 